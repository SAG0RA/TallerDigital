

module paramCalculator_tb ();


endmodule